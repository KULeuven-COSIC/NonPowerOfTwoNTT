`timescale 1ns / 1ps


module merged_permutation #(  
    parameter SIZE = 257,
    parameter WIDTH = 32
 ) (   
  input  wire  [SIZE-1:0][WIDTH-1:0] input_list,
  input  wire  [2:0]                 perm_select,
  output wire  [SIZE-1:0][WIDTH-1:0] output_list
);  
    wire [SIZE*WIDTH-1:0] permutation [0:6];
    
    assign permutation[0] = {input_list[0], input_list[256], input_list[255], input_list[254], input_list[253], input_list[252], input_list[251], input_list[250], input_list[249], input_list[248], input_list[247], input_list[246], input_list[245], input_list[244], input_list[243], input_list[242], input_list[241], input_list[240], input_list[239], input_list[238], input_list[237], input_list[236], input_list[235], input_list[234], input_list[233], input_list[232], input_list[231], input_list[230], input_list[229], input_list[228], input_list[227], input_list[226], input_list[225], input_list[224], input_list[223], input_list[222], input_list[221], input_list[220], input_list[219], input_list[218], input_list[217], input_list[216], input_list[215], input_list[214], input_list[213], input_list[212], input_list[211], input_list[210], input_list[209], input_list[208], input_list[207], input_list[206], input_list[205], input_list[204], input_list[203], input_list[202], input_list[201], input_list[200], input_list[199], input_list[198], input_list[197], input_list[196], input_list[195], input_list[194], input_list[193], input_list[192], input_list[191], input_list[190], input_list[189], input_list[188], input_list[187], input_list[186], input_list[185], input_list[184], input_list[183], input_list[182], input_list[181], input_list[180], input_list[179], input_list[178], input_list[177], input_list[176], input_list[175], input_list[174], input_list[173], input_list[172], input_list[171], input_list[170], input_list[169], input_list[168], input_list[167], input_list[166], input_list[165], input_list[164], input_list[163], input_list[162], input_list[161], input_list[160], input_list[159], input_list[158], input_list[157], input_list[156], input_list[155], input_list[154], input_list[153], input_list[152], input_list[151], input_list[150], input_list[149], input_list[148], input_list[147], input_list[146], input_list[145], input_list[144], input_list[143], input_list[142], input_list[141], input_list[140], input_list[139], input_list[138], input_list[137], input_list[136], input_list[135], input_list[134], input_list[133], input_list[132], input_list[131], input_list[130], input_list[129], input_list[128], input_list[127], input_list[126], input_list[125], input_list[124], input_list[123], input_list[122], input_list[121], input_list[120], input_list[119], input_list[118], input_list[117], input_list[116], input_list[115], input_list[114], input_list[113], input_list[112], input_list[111], input_list[110], input_list[109], input_list[108], input_list[107], input_list[106], input_list[105], input_list[104], input_list[103], input_list[102], input_list[101], input_list[100], input_list[99], input_list[98], input_list[97], input_list[96], input_list[95], input_list[94], input_list[93], input_list[92], input_list[91], input_list[90], input_list[89], input_list[88], input_list[87], input_list[86], input_list[85], input_list[84], input_list[83], input_list[82], input_list[81], input_list[80], input_list[79], input_list[78], input_list[77], input_list[76], input_list[75], input_list[74], input_list[73], input_list[72], input_list[71], input_list[70], input_list[69], input_list[68], input_list[67], input_list[66], input_list[65], input_list[64], input_list[63], input_list[62], input_list[61], input_list[60], input_list[59], input_list[58], input_list[57], input_list[56], input_list[55], input_list[54], input_list[53], input_list[52], input_list[51], input_list[50], input_list[49], input_list[48], input_list[47], input_list[46], input_list[45], input_list[44], input_list[43], input_list[42], input_list[41], input_list[40], input_list[39], input_list[38], input_list[37], input_list[36], input_list[35], input_list[34], input_list[33], input_list[32], input_list[31], input_list[30], input_list[29], input_list[28], input_list[27], input_list[26], input_list[25], input_list[24], input_list[23], input_list[22], input_list[21], input_list[20], input_list[19], input_list[18], input_list[17], input_list[16], input_list[15], input_list[14], input_list[13], input_list[12], input_list[11], input_list[10], input_list[9], input_list[8], input_list[7], input_list[6], input_list[5], input_list[4], input_list[3], input_list[2], input_list[1]};
    assign permutation[1] = {input_list[0], input_list[17], input_list[34], input_list[51], input_list[68], input_list[85], input_list[102], input_list[119], input_list[136], input_list[153], input_list[170], input_list[187], input_list[204], input_list[221], input_list[238], 64'b0, input_list[254], input_list[253], input_list[252], input_list[251], input_list[250], input_list[249], input_list[248], input_list[247], input_list[246], input_list[245], input_list[244], input_list[243], input_list[242], input_list[241], input_list[240], input_list[239], input_list[237], input_list[236], input_list[235], input_list[234], input_list[233], input_list[232], input_list[231], input_list[230], input_list[229], input_list[228], input_list[227], input_list[226], input_list[225], input_list[224], input_list[223], input_list[222], input_list[220], input_list[219], input_list[218], input_list[217], input_list[216], input_list[215], input_list[214], input_list[213], input_list[212], input_list[211], input_list[210], input_list[209], input_list[208], input_list[207], input_list[206], input_list[205], input_list[203], input_list[202], input_list[201], input_list[200], input_list[199], input_list[198], input_list[197], input_list[196], input_list[195], input_list[194], input_list[193], input_list[192], input_list[191], input_list[190], input_list[189], input_list[188], input_list[186], input_list[185], input_list[184], input_list[183], input_list[182], input_list[181], input_list[180], input_list[179], input_list[178], input_list[177], input_list[176], input_list[175], input_list[174], input_list[173], input_list[172], input_list[171], input_list[169], input_list[168], input_list[167], input_list[166], input_list[165], input_list[164], input_list[163], input_list[162], input_list[161], input_list[160], input_list[159], input_list[158], input_list[157], input_list[156], input_list[155], input_list[154], input_list[152], input_list[151], input_list[150], input_list[149], input_list[148], input_list[147], input_list[146], input_list[145], input_list[144], input_list[143], input_list[142], input_list[141], input_list[140], input_list[139], input_list[138], input_list[137], input_list[135], input_list[134], input_list[133], input_list[132], input_list[131], input_list[130], input_list[129], input_list[128], input_list[127], input_list[126], input_list[125], input_list[124], input_list[123], input_list[122], input_list[121], input_list[120], input_list[118], input_list[117], input_list[116], input_list[115], input_list[114], input_list[113], input_list[112], input_list[111], input_list[110], input_list[109], input_list[108], input_list[107], input_list[106], input_list[105], input_list[104], input_list[103], input_list[101], input_list[100], input_list[99], input_list[98], input_list[97], input_list[96], input_list[95], input_list[94], input_list[93], input_list[92], input_list[91], input_list[90], input_list[89], input_list[88], input_list[87], input_list[86], input_list[84], input_list[83], input_list[82], input_list[81], input_list[80], input_list[79], input_list[78], input_list[77], input_list[76], input_list[75], input_list[74], input_list[73], input_list[72], input_list[71], input_list[70], input_list[69], input_list[67], input_list[66], input_list[65], input_list[64], input_list[63], input_list[62], input_list[61], input_list[60], input_list[59], input_list[58], input_list[57], input_list[56], input_list[55], input_list[54], input_list[53], input_list[52], input_list[50], input_list[49], input_list[48], input_list[47], input_list[46], input_list[45], input_list[44], input_list[43], input_list[42], input_list[41], input_list[40], input_list[39], input_list[38], input_list[37], input_list[36], input_list[35], input_list[33], input_list[32], input_list[31], input_list[30], input_list[29], input_list[28], input_list[27], input_list[26], input_list[25], input_list[24], input_list[23], input_list[22], input_list[21], input_list[20], input_list[19], input_list[18], input_list[16], input_list[15], input_list[14], input_list[13], input_list[12], input_list[11], input_list[10], input_list[9], input_list[8], input_list[7], input_list[6], input_list[5], input_list[4], input_list[3], input_list[2], input_list[1]};
    assign permutation[2] = {input_list[0], input_list[5], input_list[10], input_list[15], input_list[20], input_list[25], input_list[30], input_list[35], input_list[40], input_list[45], input_list[50], input_list[55], input_list[60], input_list[65], input_list[70], input_list[75], input_list[80], input_list[85], input_list[90], input_list[95], input_list[100], input_list[105], input_list[110], input_list[115], input_list[120], input_list[125], input_list[130], input_list[135], input_list[140], input_list[145], input_list[150], input_list[155], input_list[160], input_list[165], input_list[170], input_list[175], input_list[180], input_list[185], input_list[190], input_list[195], input_list[200], input_list[205], input_list[210], input_list[215], input_list[220], input_list[225], input_list[230], input_list[235], input_list[240], input_list[245], input_list[250], 64'b0, input_list[254], input_list[253], input_list[252], input_list[251], input_list[249], input_list[248], input_list[247], input_list[246], input_list[244], input_list[243], input_list[242], input_list[241], input_list[239], input_list[238], input_list[237], input_list[236], input_list[234], input_list[233], input_list[232], input_list[231], input_list[229], input_list[228], input_list[227], input_list[226], input_list[224], input_list[223], input_list[222], input_list[221], input_list[219], input_list[218], input_list[217], input_list[216], input_list[214], input_list[213], input_list[212], input_list[211], input_list[209], input_list[208], input_list[207], input_list[206], input_list[204], input_list[203], input_list[202], input_list[201], input_list[199], input_list[198], input_list[197], input_list[196], input_list[194], input_list[193], input_list[192], input_list[191], input_list[189], input_list[188], input_list[187], input_list[186], input_list[184], input_list[183], input_list[182], input_list[181], input_list[179], input_list[178], input_list[177], input_list[176], input_list[174], input_list[173], input_list[172], input_list[171], input_list[169], input_list[168], input_list[167], input_list[166], input_list[164], input_list[163], input_list[162], input_list[161], input_list[159], input_list[158], input_list[157], input_list[156], input_list[154], input_list[153], input_list[152], input_list[151], input_list[149], input_list[148], input_list[147], input_list[146], input_list[144], input_list[143], input_list[142], input_list[141], input_list[139], input_list[138], input_list[137], input_list[136], input_list[134], input_list[133], input_list[132], input_list[131], input_list[129], input_list[128], input_list[127], input_list[126], input_list[124], input_list[123], input_list[122], input_list[121], input_list[119], input_list[118], input_list[117], input_list[116], input_list[114], input_list[113], input_list[112], input_list[111], input_list[109], input_list[108], input_list[107], input_list[106], input_list[104], input_list[103], input_list[102], input_list[101], input_list[99], input_list[98], input_list[97], input_list[96], input_list[94], input_list[93], input_list[92], input_list[91], input_list[89], input_list[88], input_list[87], input_list[86], input_list[84], input_list[83], input_list[82], input_list[81], input_list[79], input_list[78], input_list[77], input_list[76], input_list[74], input_list[73], input_list[72], input_list[71], input_list[69], input_list[68], input_list[67], input_list[66], input_list[64], input_list[63], input_list[62], input_list[61], input_list[59], input_list[58], input_list[57], input_list[56], input_list[54], input_list[53], input_list[52], input_list[51], input_list[49], input_list[48], input_list[47], input_list[46], input_list[44], input_list[43], input_list[42], input_list[41], input_list[39], input_list[38], input_list[37], input_list[36], input_list[34], input_list[33], input_list[32], input_list[31], input_list[29], input_list[28], input_list[27], input_list[26], input_list[24], input_list[23], input_list[22], input_list[21], input_list[19], input_list[18], input_list[17], input_list[16], input_list[14], input_list[13], input_list[12], input_list[11], input_list[9], input_list[8], input_list[7], input_list[6], input_list[4], input_list[3], input_list[2], input_list[1]};
    assign permutation[3] = 'hx;
    assign permutation[4] = {input_list[0], input_list[86], input_list[171], input_list[91], input_list[166], input_list[170], input_list[87], input_list[150], input_list[107], input_list[182], input_list[75], input_list[85], input_list[172], input_list[43], input_list[214], input_list[174], input_list[83], input_list[80], input_list[177], input_list[252], input_list[5], input_list[194], input_list[63], input_list[20], input_list[237], input_list[247], input_list[10], input_list[97], input_list[160], input_list[40], input_list[217], input_list[126], input_list[131], input_list[55], input_list[202], input_list[109], input_list[148], input_list[37], input_list[220], input_list[78], input_list[179], input_list[218], input_list[39], input_list[147], input_list[110], input_list[156], input_list[101], input_list[183], input_list[74], input_list[93], input_list[164], input_list[203], input_list[54], input_list[142], input_list[115], input_list[216], input_list[41], input_list[149], input_list[108], input_list[71], input_list[186], input_list[175], input_list[82], input_list[230], input_list[27], input_list[238], input_list[19], input_list[210], input_list[47], input_list[76], input_list[181], input_list[188], input_list[69], input_list[163], input_list[94], input_list[38], input_list[219], input_list[119], input_list[138], input_list[105], input_list[152], input_list[66], input_list[191], input_list[28], input_list[229], input_list[250], input_list[7], input_list[145], input_list[112], input_list[56], input_list[201], input_list[125], input_list[132], input_list[33], input_list[224], input_list[14], input_list[243], input_list[206], input_list[51], input_list[212], input_list[45], input_list[204], input_list[53], input_list[180], input_list[77], input_list[167], input_list[90], input_list[102], input_list[155], input_list[103], input_list[154], input_list[106], input_list[151], input_list[96], input_list[161], input_list[251], input_list[6], input_list[130], input_list[127], input_list[24], input_list[233], input_list[245], input_list[12], input_list[65], input_list[192], input_list[48], input_list[209], input_list[254], input_list[3], input_list[200], input_list[57], input_list[116], input_list[141], input_list[228], input_list[29], input_list[50], input_list[207], input_list[232], input_list[25], input_list[114], input_list[143], input_list[100], input_list[157], input_list[58], input_list[199], input_list[198], input_list[59], input_list[84], input_list[173], input_list[236], input_list[21], input_list[178], input_list[79], input_list[168], input_list[89], input_list[118], input_list[139], input_list[99], input_list[158], input_list[42], input_list[215], input_list[104], input_list[153], input_list[122], input_list[135], input_list[98], input_list[159], input_list[26], input_list[231], input_list[244], input_list[13], input_list[49], input_list[208], input_list[52], input_list[205], input_list[61], input_list[196], input_list[31], input_list[226], input_list[239], input_list[18], input_list[133], input_list[124], input_list[72], input_list[185], input_list[221], input_list[36], input_list[195], input_list[62], input_list[144], input_list[113], input_list[248], input_list[9], input_list[165], input_list[92], input_list[70], input_list[187], input_list[111], input_list[146], input_list[234], input_list[23], input_list[140], input_list[117], input_list[184], input_list[73], input_list[211], input_list[46], input_list[35], input_list[222], input_list[22], input_list[235], input_list[95], input_list[162], input_list[169], input_list[88], input_list[134], input_list[123], input_list[190], input_list[67], input_list[213], input_list[44], input_list[11], input_list[246], input_list[176], input_list[81], input_list[240], input_list[17], input_list[242], input_list[15], input_list[68], input_list[189], input_list[60], input_list[197], input_list[227], input_list[30], input_list[34], input_list[223], input_list[120], input_list[137], input_list[121], input_list[136], input_list[32], input_list[225], input_list[255], input_list[2], input_list[129], input_list[128], input_list[8], input_list[249], input_list[253], input_list[4], input_list[193], input_list[64], input_list[16], input_list[241], input_list[256], input_list[1]};
    assign permutation[5] = {input_list[0], input_list[51], input_list[17], input_list[68], input_list[34], input_list[85], input_list[136], input_list[102], input_list[153], input_list[119], input_list[170], input_list[221], input_list[187], input_list[238], input_list[204], 64'b0, input_list[244], input_list[249], input_list[194], input_list[214], input_list[199], input_list[209], input_list[184], input_list[224], input_list[189], input_list[219], input_list[229], input_list[179], input_list[174], input_list[234], input_list[254], input_list[239], input_list[193], input_list[198], input_list[228], input_list[248], input_list[233], input_list[243], input_list[218], input_list[173], input_list[223], input_list[253], input_list[178], input_list[213], input_list[208], input_list[183], input_list[203], input_list[188], input_list[227], input_list[232], input_list[177], input_list[197], input_list[182], input_list[192], input_list[252], input_list[207], input_list[172], input_list[202], input_list[212], input_list[247], input_list[242], input_list[217], input_list[237], input_list[222], input_list[176], input_list[181], input_list[211], input_list[231], input_list[216], input_list[226], input_list[201], input_list[241], input_list[206], input_list[236], input_list[246], input_list[196], input_list[191], input_list[251], input_list[186], input_list[171], input_list[210], input_list[215], input_list[245], input_list[180], input_list[250], input_list[175], input_list[235], input_list[190], input_list[240], input_list[185], input_list[195], input_list[230], input_list[225], input_list[200], input_list[220], input_list[205], input_list[159], input_list[164], input_list[109], input_list[129], input_list[114], input_list[124], input_list[99], input_list[139], input_list[104], input_list[134], input_list[144], input_list[94], input_list[89], input_list[149], input_list[169], input_list[154], input_list[108], input_list[113], input_list[143], input_list[163], input_list[148], input_list[158], input_list[133], input_list[88], input_list[138], input_list[168], input_list[93], input_list[128], input_list[123], input_list[98], input_list[118], input_list[103], input_list[142], input_list[147], input_list[92], input_list[112], input_list[97], input_list[107], input_list[167], input_list[122], input_list[87], input_list[117], input_list[127], input_list[162], input_list[157], input_list[132], input_list[152], input_list[137], input_list[91], input_list[96], input_list[126], input_list[146], input_list[131], input_list[141], input_list[116], input_list[156], input_list[121], input_list[151], input_list[161], input_list[111], input_list[106], input_list[166], input_list[101], input_list[86], input_list[125], input_list[130], input_list[160], input_list[95], input_list[165], input_list[90], input_list[150], input_list[105], input_list[155], input_list[100], input_list[110], input_list[145], input_list[140], input_list[115], input_list[135], input_list[120], input_list[74], input_list[79], input_list[24], input_list[44], input_list[29], input_list[39], input_list[14], input_list[54], input_list[19], input_list[49], input_list[59], input_list[9], input_list[4], input_list[64], input_list[84], input_list[69], input_list[23], input_list[28], input_list[58], input_list[78], input_list[63], input_list[73], input_list[48], input_list[3], input_list[53], input_list[83], input_list[8], input_list[43], input_list[38], input_list[13], input_list[33], input_list[18], input_list[57], input_list[62], input_list[7], input_list[27], input_list[12], input_list[22], input_list[82], input_list[37], input_list[2], input_list[32], input_list[42], input_list[77], input_list[72], input_list[47], input_list[67], input_list[52], input_list[6], input_list[11], input_list[41], input_list[61], input_list[46], input_list[56], input_list[31], input_list[71], input_list[36], input_list[66], input_list[76], input_list[26], input_list[21], input_list[81], input_list[16], input_list[1], input_list[40], input_list[45], input_list[75], input_list[10], input_list[80], input_list[5], input_list[65], input_list[20], input_list[70], input_list[15], input_list[25], input_list[60], input_list[55], input_list[30], input_list[50], input_list[35]};
    assign permutation[6] = {input_list[0], input_list[1], input_list[2], input_list[3], input_list[4], input_list[5], input_list[6], input_list[7], input_list[8], input_list[9], input_list[10], input_list[11], input_list[12], input_list[13], input_list[14], input_list[15], input_list[16], input_list[85], input_list[86], input_list[87], input_list[88], input_list[89], input_list[90], input_list[91], input_list[92], input_list[93], input_list[94], input_list[95], input_list[96], input_list[97], input_list[98], input_list[99], input_list[100], input_list[101], input_list[170], input_list[171], input_list[172], input_list[173], input_list[174], input_list[175], input_list[176], input_list[177], input_list[178], input_list[179], input_list[180], input_list[181], input_list[182], input_list[183], input_list[184], input_list[185], input_list[186], 64'b0, input_list[237], input_list[220], input_list[254], input_list[203], input_list[236], input_list[219], input_list[253], input_list[202], input_list[235], input_list[218], input_list[252], input_list[201], input_list[234], input_list[217], input_list[251], input_list[200], input_list[233], input_list[216], input_list[250], input_list[199], input_list[232], input_list[215], input_list[249], input_list[198], input_list[231], input_list[214], input_list[248], input_list[197], input_list[230], input_list[213], input_list[247], input_list[196], input_list[229], input_list[212], input_list[246], input_list[195], input_list[228], input_list[211], input_list[245], input_list[194], input_list[227], input_list[210], input_list[244], input_list[193], input_list[226], input_list[209], input_list[243], input_list[192], input_list[225], input_list[208], input_list[242], input_list[191], input_list[224], input_list[207], input_list[241], input_list[190], input_list[223], input_list[206], input_list[240], input_list[189], input_list[222], input_list[205], input_list[239], input_list[188], input_list[221], input_list[204], input_list[238], input_list[187], input_list[152], input_list[135], input_list[169], input_list[118], input_list[151], input_list[134], input_list[168], input_list[117], input_list[150], input_list[133], input_list[167], input_list[116], input_list[149], input_list[132], input_list[166], input_list[115], input_list[148], input_list[131], input_list[165], input_list[114], input_list[147], input_list[130], input_list[164], input_list[113], input_list[146], input_list[129], input_list[163], input_list[112], input_list[145], input_list[128], input_list[162], input_list[111], input_list[144], input_list[127], input_list[161], input_list[110], input_list[143], input_list[126], input_list[160], input_list[109], input_list[142], input_list[125], input_list[159], input_list[108], input_list[141], input_list[124], input_list[158], input_list[107], input_list[140], input_list[123], input_list[157], input_list[106], input_list[139], input_list[122], input_list[156], input_list[105], input_list[138], input_list[121], input_list[155], input_list[104], input_list[137], input_list[120], input_list[154], input_list[103], input_list[136], input_list[119], input_list[153], input_list[102], input_list[67], input_list[50], input_list[84], input_list[33], input_list[66], input_list[49], input_list[83], input_list[32], input_list[65], input_list[48], input_list[82], input_list[31], input_list[64], input_list[47], input_list[81], input_list[30], input_list[63], input_list[46], input_list[80], input_list[29], input_list[62], input_list[45], input_list[79], input_list[28], input_list[61], input_list[44], input_list[78], input_list[27], input_list[60], input_list[43], input_list[77], input_list[26], input_list[59], input_list[42], input_list[76], input_list[25], input_list[58], input_list[41], input_list[75], input_list[24], input_list[57], input_list[40], input_list[74], input_list[23], input_list[56], input_list[39], input_list[73], input_list[22], input_list[55], input_list[38], input_list[72], input_list[21], input_list[54], input_list[37], input_list[71], input_list[20], input_list[53], input_list[36], input_list[70], input_list[19], input_list[52], input_list[35], input_list[69], input_list[18], input_list[51], input_list[34], input_list[68], input_list[17]};

    
    assign output_list = permutation[perm_select];
         
endmodule